library verilog;
use verilog.vl_types.all;
entity sv_class_ex is
end sv_class_ex;
