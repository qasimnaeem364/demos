library verilog;
use verilog.vl_types.all;
entity top_sv_unit is
end top_sv_unit;
