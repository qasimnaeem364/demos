library verilog;
use verilog.vl_types.all;
entity usb_pkg is
end usb_pkg;
